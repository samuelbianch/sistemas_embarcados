module circuito(a, b, c, xor1, s);

	input a, b, c;
	output xor1, s;

	xor(xor1, a, b);
	and(s, xor1, c);

endmodule
