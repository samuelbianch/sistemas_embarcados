module  and_gate_2(a, b, s);

  input a, b;
  output s;
  assign s = a & b;

endmodule
