module and_gate_a(a, b, s);

	input a, b;
	output s;

	and(s, a, b);

endmodule
